`include "uvm_macros.svh"
import uvm_pkg::*;

module tb;
  initial begin
    `uvm_info("TB_TOP", "First RTL: Test_Bench_Top", UVM_MEDIUM);
  end
endmodule
